module memory

import external
import internal